* Equivalent circuit model for JWS_InductorRed_v2.ckt
.SUBCKT JWS_InductorRed_v2 po1
Vsp1 po1 p1 0
Vsr1 p1 pr1 0
Rp1 pr1 0 50
Ru1 u1 0 50
Fr1 u1 0 Vsr1 -1
Fu1 u1 0 Vsp1 -1
Ry1 y1 0 1
Gy1 p1 0 y1 0 -0.02
Rx1 x1 0 1
Fxc1_2 x1 0 Vx2 7.53325734982205
Cx1 x1 xm1 0.0144258823575351
Vx1 xm1 0 0
Gx1_1 x1 0 u1 0 -1.2406808347684
Rx2 x2 0 1
Fxc2_1 x2 0 Vx1 -0.109129748189251
Cx2 x2 xm2 0.0144258823575351
Vx2 xm2 0 0
Gx2_1 x2 0 u1 0 0.135395187081506
Rx3 x3 0 1
Cx3 x3 0 0.0545063822621616
Gx3_1 x3 0 u1 0 -2.18390144792024
Rx4 x4 0 1
Fxc4_5 x4 0 Vx5 395.931609951382
Cx4 x4 xm4 9.2663822324964e-05
Vx4 xm4 0 0
Gx4_1 x4 0 u1 0 -2.54844093535363e-05
Rx5 x5 0 1
Fxc5_4 x5 0 Vx4 -300.138552338075
Cx5 x5 xm5 9.2663822324964e-05
Vx5 xm5 0 0
Gx5_1 x5 0 u1 0 0.0076488537305613
Rx6 x6 0 1
Fxc6_7 x6 0 Vx7 4485.70686026196
Cx6 x6 xm6 8.27811924909976e-06
Vx6 xm6 0 0
Gx6_1 x6 0 u1 0 -1.6669253143261e-07
Rx7 x7 0 1
Fxc7_6 x7 0 Vx6 -3880.10266727079
Cx7 x7 xm7 8.27811924909976e-06
Vx7 xm7 0 0
Gx7_1 x7 0 u1 0 0.000646784135825789
Rx8 x8 0 1
Fxc8_9 x8 0 Vx9 2033.06944367417
Cx8 x8 xm8 1.4704310556239e-05
Vx8 xm8 0 0
Gx8_1 x8 0 u1 0 -3.84649635257523e-07
Rx9 x9 0 1
Fxc9_8 x9 0 Vx8 -3178.51479990235
Cx9 x9 xm9 1.4704310556239e-05
Vx9 xm9 0 0
Gx9_1 x9 0 u1 0 0.00122261455844308
Rx10 x10 0 1
Cx10 x10 0 6.20658031512027
Gx10_1 x10 0 u1 0 -2.03778145438967
Rx11 x11 0 1
Fxc11_12 x11 0 Vx12 403.374406351594
Cx11 x11 xm11 0.000442482271364814
Vx11 xm11 0 0
Gx11_1 x11 0 u1 0 -2.63564824163105e-05
Rx12 x12 0 1
Fxc12_11 x12 0 Vx11 -287.90190996354
Cx12 x12 xm12 0.000442482271364814
Vx12 xm12 0 0
Gx12_1 x12 0 u1 0 0.00758808162757625
Rx13 x13 0 1
Fxc13_14 x13 0 Vx14 210.374663594951
Cx13 x13 xm13 0.000177214686415986
Vx13 xm13 0 0
Gx13_1 x13 0 u1 0 -6.33916986003802e-06
Rx14 x14 0 1
Fxc14_13 x14 0 Vx13 -1171.83743906206
Cx14 x14 xm14 0.000177214686415986
Vx14 xm14 0 0
Gx14_1 x14 0 u1 0 0.00742847657456636
Rx15 x15 0 1
Fxc15_16 x15 0 Vx16 171.166055033571
Cx15 x15 xm15 9.26132475048291e-05
Vx15 xm15 0 0
Gx15_1 x15 0 u1 0 -5.19165746463756e-06
Rx16 x16 0 1
Fxc16_15 x16 0 Vx15 -1462.84612246512
Cx16 x16 xm16 9.26132475048291e-05
Vx16 xm16 0 0
Gx16_1 x16 0 u1 0 0.00759459599131213
Rx17 x17 0 1
Fxc17_18 x17 0 Vx18 328.769768578865
Cx17 x17 xm17 5.66336887557543e-05
Vx17 xm17 0 0
Gx17_1 x17 0 u1 0 -1.90348283006726e-06
Rx18 x18 0 1
Fxc18_17 x18 0 Vx17 -2278.50862110563
Cx18 x18 xm18 5.66336887557543e-05
Vx18 xm18 0 0
Gx18_1 x18 0 u1 0 0.00433710203843479
Rx19 x19 0 1
Fxc19_20 x19 0 Vx20 236.12964076412
Cx19 x19 xm19 1.22041330547248e-05
Vx19 xm19 0 0
Gx19_1 x19 0 u1 0 -8.63604142293708e-09
Rx20 x20 0 1
Fxc20_19 x20 0 Vx19 -102129.944410137
Cx20 x20 xm20 1.22041330547248e-05
Vx20 xm20 0 0
Gx20_1 x20 0 u1 0 0.000881998430448202
Gyc1_1 y1 0 x1 0 1
Gyc1_2 y1 0 x2 0 1
Gyc1_3 y1 0 x3 0 -1
Gyc1_4 y1 0 x4 0 -1
Gyc1_5 y1 0 x5 0 -1
Gyc1_6 y1 0 x6 0 -1
Gyc1_7 y1 0 x7 0 -1
Gyc1_8 y1 0 x8 0 -1
Gyc1_9 y1 0 x9 0 -1
Gyc1_10 y1 0 x10 0 1
Gyc1_11 y1 0 x11 0 1
Gyc1_12 y1 0 x12 0 -1
Gyc1_13 y1 0 x13 0 1
Gyc1_14 y1 0 x14 0 -1
Gyc1_15 y1 0 x15 0 -1
Gyc1_16 y1 0 x16 0 -1
Gyc1_17 y1 0 x17 0 -1
Gyc1_18 y1 0 x18 0 -1
Gyc1_19 y1 0 x19 0 -1
Gyc1_20 y1 0 x20 0 -1
.ENDS
