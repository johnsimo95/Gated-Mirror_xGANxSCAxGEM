* Equivalent circuit model for JWS_InductorRed_v4.ckt
.SUBCKT JWS_InductorRed_v4 po1
Vsp1 po1 p1 0
Vsr1 p1 pr1 0
Rp1 pr1 0 50
Ru1 u1 0 50
Fr1 u1 0 Vsr1 -1
Fu1 u1 0 Vsp1 -1
Ry1 y1 0 1
Gy1 p1 0 y1 0 -0.02
Rx1 x1 0 1
Fxc1_2 x1 0 Vx2 22.8080658661197
Cx1 x1 xm1 0.00332760005868646
Vx1 xm1 0 0
Gx1_1 x1 0 u1 0 -0.0150258224128132
Rx2 x2 0 1
Fxc2_1 x2 0 Vx1 -1.82399505228824
Cx2 x2 xm2 0.00332760005868646
Vx2 xm2 0 0
Gx2_1 x2 0 u1 0 0.0274070257375331
Rx3 x3 0 1
Fxc3_4 x3 0 Vx4 0.00283977501896124
Cx3 x3 xm3 0.0290921102470382
Vx3 xm3 0 0
Gx3_1 x3 0 u1 0 -1.74676983906461
Rx4 x4 0 1
Fxc4_3 x4 0 Vx3 -1.54085603773246
Cx4 x4 xm4 0.0290921102470382
Vx4 xm4 0 0
Gx4_1 x4 0 u1 0 2.69152085305167
Gyc1_1 y1 0 x1 0 -1
Gyc1_2 y1 0 x2 0 1
Gyc1_3 y1 0 x3 0 1
Gyc1_4 y1 0 x4 0 1
.ENDS
