* Equivalent circuit model for 200727_testNetworkJS_v1.ckt
.SUBCKT 200727_testNetworkJS_v1 po1
Vsp1 po1 p1 0
Vsr1 p1 pr1 0
Rp1 pr1 0 50
Ru1 u1 0 50
Fr1 u1 0 Vsr1 -1
Fu1 u1 0 Vsp1 -1
Ry1 y1 0 1
Gy1 p1 0 y1 0 -0.02
Rx1 x1 0 1
Cx1 x1 0 8.44207088386674e-12
Gx1_1 x1 0 u1 0 -1.51289136612221
Rx2 x2 0 1
Fxc2_3 x2 0 Vx3 8.00726759604801
Cx2 x2 xm2 1.11813894959864e-12
Vx2 xm2 0 0
Gx2_1 x2 0 u1 0 -0.00820706818248792
Rx3 x3 0 1
Fxc3_2 x3 0 Vx2 -20.5862823965657
Cx3 x3 xm3 1.11813894959864e-12
Vx3 xm3 0 0
Gx3_1 x3 0 u1 0 0.168953023252566
Rx4 x4 0 1
Fxc4_5 x4 0 Vx5 107.795476201096
Cx4 x4 xm4 4.71772312948075e-13
Vx4 xm4 0 0
Gx4_1 x4 0 u1 0 -0.00335916450652818
Rx5 x5 0 1
Fxc5_4 x5 0 Vx4 -13.1954111811137
Cx5 x5 xm5 4.71772312948075e-13
Vx5 xm5 0 0
Gx5_1 x5 0 u1 0 0.0443255568886423
Rx6 x6 0 1
Fxc6_7 x6 0 Vx7 2.81029851423148
Cx6 x6 xm6 5.04562498515061e-14
Vx6 xm6 0 0
Gx6_1 x6 0 u1 0 -2.75988214299181e-07
Rx7 x7 0 1
Fxc7_6 x7 0 Vx6 -46053.064025524
Cx7 x7 xm7 5.0456249851506e-14
Vx7 xm7 0 0
Gx7_1 x7 0 u1 0 0.0127101029034102
Rx8 x8 0 1
Fxc8_9 x8 0 Vx9 17749.7487987464
Cx8 x8 xm8 1.82330521684262e-14
Vx8 xm8 0 0
Gx8_1 x8 0 u1 0 -3.39640752468932e-06
Rx9 x9 0 1
Fxc9_8 x9 0 Vx8 -65.3188429155793
Cx9 x9 xm9 1.82330521684262e-14
Vx9 xm9 0 0
Gx9_1 x9 0 u1 0 0.000221849409582473
Rx10 x10 0 1
Cx10 x10 0 5.97310646437398e-10
Gx10_1 x10 0 u1 0 -2.2434998574718
Rx11 x11 0 1
Fxc11_12 x11 0 Vx12 494.599263490855
Cx11 x11 xm11 2.12403439310865e-13
Vx11 xm11 0 0
Gx11_1 x11 0 u1 0 -6.86891322290552e-08
Rx12 x12 0 1
Fxc12_11 x12 0 Vx11 -606.550897317283
Cx12 x12 xm12 2.12403439310865e-13
Vx12 xm12 0 0
Gx12_1 x12 0 u1 0 4.16634547894789e-05
Rx13 x13 0 1
Fxc13_14 x13 0 Vx14 1347.89407706854
Cx13 x13 xm13 4.35737999254938e-14
Vx13 xm13 0 0
Gx13_1 x13 0 u1 0 -1.95246466279752e-06
Rx14 x14 0 1
Fxc14_13 x14 0 Vx13 -1130.2222575025
Cx14 x14 xm14 4.35737999254937e-14
Vx14 xm14 0 0
Gx14_1 x14 0 u1 0 0.00220671901888087
Rx15 x15 0 1
Fxc15_16 x15 0 Vx16 3.56880171859102
Cx15 x15 xm15 5.46819085120128e-12
Vx15 xm15 0 0
Gx15_1 x15 0 u1 0 -0.0308303615524686
Rx16 x16 0 1
Fxc16_15 x16 0 Vx15 -20.3078765590217
Cx16 x16 xm16 5.46819085120128e-12
Vx16 xm16 0 0
Gx16_1 x16 0 u1 0 0.62609917667754
Rx17 x17 0 1
Fxc17_18 x17 0 Vx18 9.82687829820278
Cx17 x17 xm17 8.28540469734822e-12
Vx17 xm17 0 0
Gx17_1 x17 0 u1 0 -0.388389633111233
Rx18 x18 0 1
Fxc18_17 x18 0 Vx17 -1.51388199113502
Cx18 x18 xm18 8.28540469734822e-12
Vx18 xm18 0 0
Gx18_1 x18 0 u1 0 0.587976071110635
Rx19 x19 0 1
Fxc19_20 x19 0 Vx20 2445.75323044656
Cx19 x19 xm19 7.31288393807337e-15
Vx19 xm19 0 0
Gx19_1 x19 0 u1 0 -2.55578195983261e-07
Rx20 x20 0 1
Fxc20_19 x20 0 Vx19 -4227.87296058262
Cx20 x20 xm20 7.31288393807337e-15
Vx20 xm20 0 0
Gx20_1 x20 0 u1 0 0.00108055214411212
Rx21 x21 0 1
Fxc21_22 x21 0 Vx22 3969.90930100717
Cx21 x21 xm21 3.43169342932507e-15
Vx21 xm21 0 0
Gx21_1 x21 0 u1 0 -3.10247465268833e-08
Rx22 x22 0 1
Fxc22_21 x22 0 Vx21 -12396.8871452701
Cx22 x22 xm22 3.43169342932507e-15
Vx22 xm22 0 0
Gx22_1 x22 0 u1 0 0.000384610281404383
Rx23 x23 0 1
Fxc23_24 x23 0 Vx24 803.598631995011
Cx23 x23 xm23 8.83713688313861e-15
Vx23 xm23 0 0
Gx23_1 x23 0 u1 0 -1.1039323319929e-07
Rx24 x24 0 1
Fxc24_23 x24 0 Vx23 -10511.4611731532
Cx24 x24 xm24 8.83713688313861e-15
Vx24 xm24 0 0
Gx24_1 x24 0 u1 0 0.00116039418455318
Gyc1_1 y1 0 x1 0 1
Gyc1_2 y1 0 x2 0 -1
Gyc1_3 y1 0 x3 0 -1
Gyc1_4 y1 0 x4 0 -1
Gyc1_5 y1 0 x5 0 -1
Gyc1_6 y1 0 x6 0 1
Gyc1_7 y1 0 x7 0 1
Gyc1_8 y1 0 x8 0 -1
Gyc1_9 y1 0 x9 0 1
Gyc1_10 y1 0 x10 0 -1
Gyc1_11 y1 0 x11 0 -1
Gyc1_12 y1 0 x12 0 1
Gyc1_13 y1 0 x13 0 1
Gyc1_14 y1 0 x14 0 1
Gyc1_15 y1 0 x15 0 -1
Gyc1_16 y1 0 x16 0 1
Gyc1_17 y1 0 x17 0 -1
Gyc1_18 y1 0 x18 0 -1
Gyc1_19 y1 0 x19 0 -1
Gyc1_20 y1 0 x20 0 -1
Gyc1_21 y1 0 x21 0 -1
Gyc1_22 y1 0 x22 0 -1
Gyc1_23 y1 0 x23 0 -1
Gyc1_24 y1 0 x24 0 -1
.ENDS
