* Equivalent circuit model for testNetworkJS_v6.ckt
.SUBCKT testNetworkJS_v6 po1
Vsp1 po1 p1 0
Vsr1 p1 pr1 0
Rp1 pr1 0 50
Ru1 u1 0 50
Fr1 u1 0 Vsr1 -1
Fu1 u1 0 Vsp1 -1
Ry1 y1 0 1
Gy1 p1 0 y1 0 -0.02
Rx1 x1 0 1
Fxc1_2 x1 0 Vx2 153184923.364426
Cx1 x1 xm1 6.27732293704952e-16
Vx1 xm1 0 0
Gx1_1 x1 0 u1 0 -0.000623992976817302
Rx2 x2 0 1
Fxc2_1 x2 0 Vx1 -2.6206901031631
Cx2 x2 xm2 6.27732293704952e-16
Vx2 xm2 0 0
Gx2_1 x2 0 u1 0 0.00163529221878838
Rx3 x3 0 1
Fxc3_4 x3 0 Vx4 4689812316488.47
Cx3 x3 xm3 3.66203687247383e-19
Vx3 xm3 0 0
Gx3_1 x3 0 u1 0 -4.87109075524666e-08
Rx4 x4 0 1
Fxc4_3 x4 0 Vx3 -498.62574945995
Cx4 x4 xm4 3.66203687247383e-19
Vx4 xm4 0 0
Gx4_1 x4 0 u1 0 2.4288512785223e-05
Rx5 x5 0 1
Fxc5_6 x5 0 Vx6 647069123097.662
Cx5 x5 xm5 1.32056042554838e-18
Vx5 xm5 0 0
Gx5_1 x5 0 u1 0 -3.34233127687062e-08
Rx6 x6 0 1
Fxc6_5 x6 0 Vx5 -293.257176232599
Cx6 x6 xm6 1.32056042554838e-18
Vx6 xm6 0 0
Gx6_1 x6 0 u1 0 9.80162632288974e-06
Rx7 x7 0 1
Fxc7_8 x7 0 Vx8 443305410569.563
Cx7 x7 xm7 1.05583730024997e-18
Vx7 xm7 0 0
Gx7_1 x7 0 u1 0 -6.30598622339785e-09
Rx8 x8 0 1
Fxc8_7 x8 0 Vx7 -779.582240962369
Cx8 x8 xm8 1.05583730024997e-18
Vx8 xm8 0 0
Gx8_1 x8 0 u1 0 4.91603487151432e-06
Rx9 x9 0 1
Fxc9_10 x9 0 Vx10 3048980740.55967
Cx9 x9 xm9 3.74619055735731e-16
Vx9 xm9 0 0
Gx9_1 x9 0 u1 0 -0.000103065248906228
Rx10 x10 0 1
Fxc10_9 x10 0 Vx9 -5.95012583779279
Cx10 x10 xm10 3.74619055735731e-16
Vx10 xm10 0 0
Gx10_1 x10 0 u1 0 0.000613251200495492
Rx11 x11 0 1
Fxc11_12 x11 0 Vx12 204937826314.78
Cx11 x11 xm11 1.16496576106882e-18
Vx11 xm11 0 0
Gx11_1 x11 0 u1 0 -2.63451909058408e-09
Rx12 x12 0 1
Fxc12_11 x12 0 Vx11 -2370.99223467072
Cx12 x12 xm12 1.16496576106882e-18
Vx12 xm12 0 0
Gx12_1 x12 0 u1 0 6.24642430586662e-06
Rx13 x13 0 1
Fxc13_14 x13 0 Vx14 96400216283349
Cx13 x13 xm13 1.21879493375187e-18
Vx13 xm13 0 0
Gx13_1 x13 0 u1 0 -7.4894115587095e-07
Rx14 x14 0 1
Fxc14_13 x14 0 Vx13 -7.18763411831909
Cx14 x14 xm14 1.21879493375187e-18
Vx14 xm14 0 0
Gx14_1 x14 0 u1 0 5.38311500455137e-06
Rx15 x15 0 1
Fxc15_16 x15 0 Vx16 146669700408.168
Cx15 x15 xm15 1.69527587992011e-17
Vx15 xm15 0 0
Gx15_1 x15 0 u1 0 -1.64519304738761e-07
Rx16 x16 0 1
Fxc16_15 x16 0 Vx15 -21.8791108493224
Cx16 x16 xm16 1.69527587992011e-17
Vx16 xm16 0 0
Gx16_1 x16 0 u1 0 3.59953610523282e-06
Gyc1_1 y1 0 x1 0 -1
Gyc1_2 y1 0 x2 0 -1
Gyc1_3 y1 0 x3 0 -1
Gyc1_4 y1 0 x4 0 1
Gyc1_5 y1 0 x5 0 -1
Gyc1_6 y1 0 x6 0 1
Gyc1_7 y1 0 x7 0 -1
Gyc1_8 y1 0 x8 0 -1
Gyc1_9 y1 0 x9 0 -1
Gyc1_10 y1 0 x10 0 1
Gyc1_11 y1 0 x11 0 -1
Gyc1_12 y1 0 x12 0 1
Gyc1_13 y1 0 x13 0 -1
Gyc1_14 y1 0 x14 0 1
Gyc1_15 y1 0 x15 0 -1
Gyc1_16 y1 0 x16 0 -1
.ENDS
