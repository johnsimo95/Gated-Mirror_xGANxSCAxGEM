* Equivalent circuit model for testNetworkJS.ckt
.SUBCKT testNetworkJS po1
Vsp1 po1 p1 0
Vsr1 p1 pr1 0
Rp1 pr1 0 50
Ru1 u1 0 50
Fr1 u1 0 Vsr1 -1
Fu1 u1 0 Vsp1 -1
Ry1 y1 0 1
Gy1 p1 0 y1 0 -0.02
Rx1 x1 0 1
Fxc1_2 x1 0 Vx2 5842310400.25508
Cx1 x1 xm1 3.60252966262071e-16
Vx1 xm1 0 0
Gx1_1 x1 0 u1 0 -0.000387936275718842
Rx2 x2 0 1
Fxc2_1 x2 0 Vx1 -1.12509522261257
Cx2 x2 xm2 3.60252966262071e-16
Vx2 xm2 0 0
Gx2_1 x2 0 u1 0 0.000436465250489383
Rx3 x3 0 1
Fxc3_4 x3 0 Vx4 89375869052222.1
Cx3 x3 xm3 2.51608510162583e-18
Vx3 xm3 0 0
Gx3_1 x3 0 u1 0 -6.53307527035151e-07
Rx4 x4 0 1
Fxc4_3 x4 0 Vx3 -4.49965724638967
Cx4 x4 xm4 2.51608510162583e-18
Vx4 xm4 0 0
Gx4_1 x4 0 u1 0 2.93965994814463e-06
Rx5 x5 0 1
Fxc5_6 x5 0 Vx6 375489836119025
Cx5 x5 xm5 2.45170974945349e-19
Vx5 xm5 0 0
Gx5_1 x5 0 u1 0 -2.63486792791916e-09
Rx6 x6 0 1
Fxc6_5 x6 0 Vx5 -128.678674984654
Cx6 x6 xm6 2.45170974945349e-19
Vx6 xm6 0 0
Gx6_1 x6 0 u1 0 3.39051313724198e-07
Rx7 x7 0 1
Cx7 x7 0 31.627559508263
Gx7_1 x7 0 u1 0 -2497168173054.67
Gyc1_1 y1 0 x1 0 -1
Gyc1_2 y1 0 x2 0 -1
Gyc1_3 y1 0 x3 0 -1
Gyc1_4 y1 0 x4 0 -1
Gyc1_5 y1 0 x5 0 -1
Gyc1_6 y1 0 x6 0 1
Gyc1_7 y1 0 x7 0 -1
.ENDS
