* Equivalent circuit model for testNetworkJS_v6.ckt
.SUBCKT testNetworkJS_v6 po1
Vsp1 po1 p1 0
Vsr1 p1 pr1 0
Rp1 pr1 0 50
Ru1 u1 0 50
Fr1 u1 0 Vsr1 -1
Fu1 u1 0 Vsp1 -1
Ry1 y1 0 1
Gy1 p1 0 y1 0 -0.02
Rx1 x1 0 1
Fxc1_2 x1 0 Vx2 875270363.357462
Cx1 x1 xm1 2.8780110388541e-16
Vx1 xm1 0 0
Gx1_1 x1 0 u1 0 -0.000506667242172905
Rx2 x2 0 1
Fxc2_1 x2 0 Vx1 -1.68351187559024
Cx2 x2 xm2 2.8780110388541e-16
Vx2 xm2 0 0
Gx2_1 x2 0 u1 0 0.000852980319170643
Rx3 x3 0 1
Fxc3_4 x3 0 Vx4 161742262338743
Cx3 x3 xm3 5.63016379415366e-20
Vx3 xm3 0 0
Gx3_1 x3 0 u1 0 -7.43634769151773e-09
Rx4 x4 0 1
Fxc4_3 x4 0 Vx3 -611.645880019828
Cx4 x4 xm4 5.63016379415366e-20
Vx4 xm4 0 0
Gx4_1 x4 0 u1 0 4.54841142791178e-06
Rx5 x5 0 1
Fxc5_6 x5 0 Vx6 545699971134.142
Cx5 x5 xm5 5.04503480463122e-18
Vx5 xm5 0 0
Gx5_1 x5 0 u1 0 -1.26201685027527e-07
Rx6 x6 0 1
Fxc6_5 x6 0 Vx5 -23.822162310129
Cx6 x6 xm6 5.04503480463122e-18
Vx6 xm6 0 0
Gx6_1 x6 0 u1 0 3.00639702453752e-06
Rx7 x7 0 1
Fxc7_8 x7 0 Vx8 8994084140.45307
Cx7 x7 xm7 6.89575256459782e-18
Vx7 xm7 0 0
Gx7_1 x7 0 u1 0 -4.07373767150656e-08
Rx8 x8 0 1
Fxc8_7 x8 0 Vx7 -900.804032622627
Cx8 x8 xm8 6.89575256459782e-18
Vx8 xm8 0 0
Gx8_1 x8 0 u1 0 3.66963932233982e-05
Rx9 x9 0 1
Fxc9_10 x9 0 Vx10 183597051.558922
Cx9 x9 xm9 4.52064952109576e-17
Vx9 xm9 0 0
Gx9_1 x9 0 u1 0 -1.58357618708977e-07
Rx10 x10 0 1
Fxc10_9 x10 0 Vx9 -1758.25105297457
Cx10 x10 xm10 4.52064952109576e-17
Vx10 xm10 0 0
Gx10_1 x10 0 u1 0 0.000278432449841604
Rx11 x11 0 1
Fxc11_12 x11 0 Vx12 95524500772607.4
Cx11 x11 xm11 9.83055925976201e-19
Vx11 xm11 0 0
Gx11_1 x11 0 u1 0 -6.05165990149426e-07
Rx12 x12 0 1
Fxc12_11 x12 0 Vx11 -11.1503120992087
Cx12 x12 xm12 9.83055925976201e-19
Vx12 xm12 0 0
Gx12_1 x12 0 u1 0 6.74778966199274e-06
Rx13 x13 0 1
Fxc13_14 x13 0 Vx14 115194894607870
Cx13 x13 xm13 2.51060190407615e-18
Vx13 xm13 0 0
Gx13_1 x13 0 u1 0 -6.51895858773719e-07
Rx14 x14 0 1
Fxc14_13 x14 0 Vx13 -3.50640123937657
Cx14 x14 xm14 2.51060190407615e-18
Vx14 xm14 0 0
Gx14_1 x14 0 u1 0 2.28580844714862e-06
Rx15 x15 0 1
Fxc15_16 x15 0 Vx16 188224115693802
Cx15 x15 xm15 1.33678494536307e-19
Vx15 xm15 0 0
Gx15_1 x15 0 u1 0 -1.43518258089593e-09
Rx16 x16 0 1
Fxc16_15 x16 0 Vx15 -863.471995820588
Cx16 x16 xm16 1.33678494536307e-19
Vx16 xm16 0 0
Gx16_1 x16 0 u1 0 1.23923996749315e-06
Rx17 x17 0 1
Cx17 x17 0 0.000639727671326046
Gx17_1 x17 0 u1 0 -50499139.2615005
Gyc1_1 y1 0 x1 0 -1
Gyc1_2 y1 0 x2 0 -1
Gyc1_3 y1 0 x3 0 -1
Gyc1_4 y1 0 x4 0 -1
Gyc1_5 y1 0 x5 0 -1
Gyc1_6 y1 0 x6 0 1
Gyc1_7 y1 0 x7 0 -1
Gyc1_8 y1 0 x8 0 -1
Gyc1_9 y1 0 x9 0 -1
Gyc1_10 y1 0 x10 0 1
Gyc1_11 y1 0 x11 0 -1
Gyc1_12 y1 0 x12 0 1
Gyc1_13 y1 0 x13 0 -1
Gyc1_14 y1 0 x14 0 -1
Gyc1_15 y1 0 x15 0 -1
Gyc1_16 y1 0 x16 0 1
Gyc1_17 y1 0 x17 0 -1
.ENDS
