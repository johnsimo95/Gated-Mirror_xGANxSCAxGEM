* Equivalent circuit model for JWS_TestNetwork_v0.ckt
.SUBCKT JWS_TestNetwork_v0 po1
Vsp1 po1 p1 0
Vsr1 p1 pr1 0
Rp1 pr1 0 50
Ru1 u1 0 50
Fr1 u1 0 Vsr1 -1
Fu1 u1 0 Vsp1 -1
Ry1 y1 0 1
Gy1 p1 0 y1 0 -0.02
Rx1 x1 0 1
Fxc1_2 x1 0 Vx2 1.49441236417188
Cx1 x1 xm1 7.62350194843161e-12
Vx1 xm1 0 0
Gx1_1 x1 0 u1 0 -0.797999729658869
Rx2 x2 0 1
Fxc2_1 x2 0 Vx1 -1.0304615403882
Cx2 x2 xm2 7.62350194843161e-12
Vx2 xm2 0 0
Gx2_1 x2 0 u1 0 0.822308030653646
Rx3 x3 0 1
Fxc3_4 x3 0 Vx4 134.972242444069
Cx3 x3 xm3 5.05165792853174e-13
Vx3 xm3 0 0
Gx3_1 x3 0 u1 0 -0.0040759360675756
Rx4 x4 0 1
Fxc4_3 x4 0 Vx3 -7.73813585498228
Cx4 x4 xm4 5.05165792853174e-13
Vx4 xm4 0 0
Gx4_1 x4 0 u1 0 0.0315401470271222
Rx5 x5 0 1
Fxc5_6 x5 0 Vx6 1749.2233852846
Cx5 x5 xm5 1.97882475535774e-14
Vx5 xm5 0 0
Gx5_1 x5 0 u1 0 -4.63882905803646e-06
Rx6 x6 0 1
Fxc6_5 x6 0 Vx5 -446.924149940254
Cx6 x6 xm6 1.97882475535774e-14
Vx6 xm6 0 0
Gx6_1 x6 0 u1 0 0.0020732047334811
Rx7 x7 0 1
Fxc7_8 x7 0 Vx8 14219.912642668
Cx7 x7 xm7 5.88311971947721e-15
Vx7 xm7 0 0
Gx7_1 x7 0 u1 0 -3.70264527454175e-07
Rx8 x8 0 1
Fxc8_7 x8 0 Vx7 -736.844586982994
Cx8 x8 xm8 5.88311971947721e-15
Vx8 xm8 0 0
Gx8_1 x8 0 u1 0 0.000272827412806425
Rx9 x9 0 1
Fxc9_10 x9 0 Vx10 193845.68638419
Cx9 x9 xm9 2.08054362171665e-16
Vx9 xm9 0 0
Gx9_1 x9 0 u1 0 -4.55678296903021e-10
Rx10 x10 0 1
Fxc10_9 x10 0 Vx9 -47519.0209906086
Cx10 x10 xm10 2.08054362171665e-16
Vx10 xm10 0 0
Gx10_1 x10 0 u1 0 2.16533865554994e-05
Rx11 x11 0 1
Cx11 x11 0 3.38196819550669e-10
Gx11_1 x11 0 u1 0 -2.41038903327483
Rx12 x12 0 1
Fxc12_13 x12 0 Vx13 15.1484946156722
Cx12 x12 xm12 9.31993415098209e-12
Vx12 xm12 0 0
Gx12_1 x12 0 u1 0 -0.264518654161207
Rx13 x13 0 1
Fxc13_12 x13 0 Vx12 -1.35664974788445
Cx13 x13 xm13 9.31993415098209e-12
Vx13 xm13 0 0
Gx13_1 x13 0 u1 0 0.358859165478537
Rx14 x14 0 1
Fxc14_15 x14 0 Vx15 5394.5426304348
Cx14 x14 xm14 2.17606443767413e-14
Vx14 xm14 0 0
Gx14_1 x14 0 u1 0 -9.22704935162211e-07
Rx15 x15 0 1
Fxc15_14 x15 0 Vx14 -768.471639526858
Cx15 x15 xm15 2.17606443767413e-14
Vx15 xm15 0 0
Gx15_1 x15 0 u1 0 0.000709072574323628
Rx16 x16 0 1
Fxc16_17 x16 0 Vx17 151368.044729615
Cx16 x16 xm16 7.90474378744846e-17
Vx16 xm16 0 0
Gx16_1 x16 0 u1 0 -1.42394011397418e-10
Rx17 x17 0 1
Fxc17_16 x17 0 Vx16 -620654.163345747
Cx17 x17 xm17 7.90474378744846e-17
Vx17 xm17 0 0
Gx17_1 x17 0 u1 0 8.83774360093092e-05
Rx18 x18 0 1
Fxc18_19 x18 0 Vx19 9.86585416165892
Cx18 x18 xm18 3.97851304101635e-12
Vx18 xm18 0 0
Gx18_1 x18 0 u1 0 -0.102687069463393
Rx19 x19 0 1
Fxc19_18 x19 0 Vx18 -4.70868205307426
Cx19 x19 xm19 3.97851304101635e-12
Vx19 xm19 0 0
Gx19_1 x19 0 u1 0 0.48352076106507
Rx20 x20 0 1
Fxc20_21 x20 0 Vx21 7308.51989794072
Cx20 x20 xm20 2.33773915563696e-15
Vx20 xm20 0 0
Gx20_1 x20 0 u1 0 -6.01662952250095e-09
Rx21 x21 0 1
Fxc21_20 x21 0 Vx20 -20311.8915897218
Cx21 x21 xm21 2.33773915563696e-15
Vx21 xm21 0 0
Gx21_1 x21 0 u1 0 0.000122209126596559
Gyc1_1 y1 0 x1 0 1
Gyc1_2 y1 0 x2 0 -1
Gyc1_3 y1 0 x3 0 -1
Gyc1_4 y1 0 x4 0 -1
Gyc1_5 y1 0 x5 0 -1
Gyc1_6 y1 0 x6 0 1
Gyc1_7 y1 0 x7 0 -1
Gyc1_8 y1 0 x8 0 -1
Gyc1_9 y1 0 x9 0 -1
Gyc1_10 y1 0 x10 0 -1
Gyc1_11 y1 0 x11 0 -1
Gyc1_12 y1 0 x12 0 -1
Gyc1_13 y1 0 x13 0 1
Gyc1_14 y1 0 x14 0 1
Gyc1_15 y1 0 x15 0 -1
Gyc1_16 y1 0 x16 0 1
Gyc1_17 y1 0 x17 0 -1
Gyc1_18 y1 0 x18 0 -1
Gyc1_19 y1 0 x19 0 -1
Gyc1_20 y1 0 x20 0 1
Gyc1_21 y1 0 x21 0 1
.ENDS
