* Equivalent circuit model for testNetworkJS_v5.ckt
.SUBCKT testNetworkJS_v5 po1
Vsp1 po1 p1 0
Vsr1 p1 pr1 0
Rp1 pr1 0 50
Ru1 u1 0 50
Fr1 u1 0 Vsr1 -1
Fu1 u1 0 Vsp1 -1
Ry1 y1 0 1
Gy1 p1 0 y1 0 -0.02
Rx1 x1 0 1
Fxc1_2 x1 0 Vx2 46006251038436.1
Cx1 x1 xm1 3.66538676574973e-18
Vx1 xm1 0 0
Gx1_1 x1 0 u1 0 -3.94556159888094e-06
Rx2 x2 0 1
Fxc2_1 x2 0 Vx1 -1.38057692502387
Cx2 x2 xm2 3.66538676574973e-18
Vx2 xm2 0 0
Gx2_1 x2 0 u1 0 5.44715129967532e-06
Rx3 x3 0 1
Fxc3_4 x3 0 Vx4 111253630881130
Cx3 x3 xm3 2.51164389003836e-18
Vx3 xm3 0 0
Gx3_1 x3 0 u1 0 -6.52154543552717e-07
Rx4 x4 0 1
Fxc4_3 x4 0 Vx3 -3.62760541805167
Cx4 x4 xm4 2.51164389003836e-18
Vx4 xm4 0 0
Gx4_1 x4 0 u1 0 2.36575935559885e-06
Rx5 x5 0 1
Fxc5_6 x5 0 Vx6 202096782264228
Cx5 x5 xm5 1.63607338792164e-19
Vx5 xm5 0 0
Gx5_1 x5 0 u1 0 -1.75833041509844e-09
Rx6 x6 0 1
Fxc6_5 x6 0 Vx5 -536.880819619885
Cx6 x6 xm6 1.63607338792164e-19
Vx6 xm6 0 0
Gx6_1 x6 0 u1 0 9.44013874420621e-07
Rx7 x7 0 1
Cx7 x7 0 0.000642452964926869
Gx7_1 x7 0 u1 0 -50726851.055196
Gyc1_1 y1 0 x1 0 -1
Gyc1_2 y1 0 x2 0 -1
Gyc1_3 y1 0 x3 0 -1
Gyc1_4 y1 0 x4 0 -1
Gyc1_5 y1 0 x5 0 -1
Gyc1_6 y1 0 x6 0 1
Gyc1_7 y1 0 x7 0 -1
.ENDS
