* Equivalent circuit model for JWS_InductorRed_v8.ckt
.SUBCKT JWS_InductorRed_v8 po1
Vsp1 po1 p1 0
Vsr1 p1 pr1 0
Rp1 pr1 0 50
Ru1 u1 0 50
Fr1 u1 0 Vsr1 -1
Fu1 u1 0 Vsp1 -1
Ry1 y1 0 1
Gy1 p1 0 y1 0 -0.02
Rx1 x1 0 1
Fxc1_2 x1 0 Vx2 7.53325734982112
Cx1 x1 xm1 1.44258823575353e-11
Vx1 xm1 0 0
Gx1_1 x1 0 u1 0 -1.24068083476842
Rx2 x2 0 1
Fxc2_1 x2 0 Vx1 -0.109129748189262
Cx2 x2 xm2 1.44258823575353e-11
Vx2 xm2 0 0
Gx2_1 x2 0 u1 0 0.135395187081521
Rx3 x3 0 1
Cx3 x3 0 5.45063822621615e-11
Gx3_1 x3 0 u1 0 -2.18390144792024
Rx4 x4 0 1
Fxc4_5 x4 0 Vx5 395.931609951365
Cx4 x4 xm4 9.26638223249673e-14
Vx4 xm4 0 0
Gx4_1 x4 0 u1 0 -2.54844093535375e-05
Rx5 x5 0 1
Fxc5_4 x5 0 Vx4 -300.138552338067
Cx5 x5 xm5 9.26638223249673e-14
Vx5 xm5 0 0
Gx5_1 x5 0 u1 0 0.00764885373056145
Rx6 x6 0 1
Fxc6_7 x6 0 Vx7 4485.70686026948
Cx6 x6 xm6 8.27811924909505e-15
Vx6 xm6 0 0
Gx6_1 x6 0 u1 0 -1.66692531432387e-07
Rx7 x7 0 1
Fxc7_6 x7 0 Vx6 -3880.1026672687
Cx7 x7 xm7 8.27811924909505e-15
Vx7 xm7 0 0
Gx7_1 x7 0 u1 0 0.000646784135824575
Rx8 x8 0 1
Fxc8_9 x8 0 Vx9 2033.06944367303
Cx8 x8 xm8 1.4704310556237e-14
Vx8 xm8 0 0
Gx8_1 x8 0 u1 0 -3.84649635257425e-07
Rx9 x9 0 1
Fxc9_8 x9 0 Vx8 -3178.51479990501
Cx9 x9 xm9 1.4704310556237e-14
Vx9 xm9 0 0
Gx9_1 x9 0 u1 0 0.00122261455844379
Rx10 x10 0 1
Cx10 x10 0 6.20658031512022e-09
Gx10_1 x10 0 u1 0 -2.03778145438966
Rx11 x11 0 1
Fxc11_12 x11 0 Vx12 403.3744063515
Cx11 x11 xm11 4.42482271364829e-13
Vx11 xm11 0 0
Gx11_1 x11 0 u1 0 -2.63564824163084e-05
Rx12 x12 0 1
Fxc12_11 x12 0 Vx11 -287.901909963588
Cx12 x12 xm12 4.42482271364829e-13
Vx12 xm12 0 0
Gx12_1 x12 0 u1 0 0.00758808162757691
Rx13 x13 0 1
Fxc13_14 x13 0 Vx14 210.374663594758
Cx13 x13 xm13 1.77214686415988e-13
Vx13 xm13 0 0
Gx13_1 x13 0 u1 0 -6.33916986003269e-06
Rx14 x14 0 1
Fxc14_13 x14 0 Vx13 -1171.83743906311
Cx14 x14 xm14 1.77214686415988e-13
Vx14 xm14 0 0
Gx14_1 x14 0 u1 0 0.00742847657456675
Rx15 x15 0 1
Fxc15_16 x15 0 Vx16 236.129640764019
Cx15 x15 xm15 1.22041330547165e-14
Vx15 xm15 0 0
Gx15_1 x15 0 u1 0 -8.63604142292239e-09
Rx16 x16 0 1
Fxc16_15 x16 0 Vx15 -102129.94441032
Cx16 x16 xm16 1.22041330547165e-14
Vx16 xm16 0 0
Gx16_1 x16 0 u1 0 0.000881998430448286
Rx17 x17 0 1
Fxc17_18 x17 0 Vx18 171.166055033454
Cx17 x17 xm17 9.26132475048371e-14
Vx17 xm17 0 0
Gx17_1 x17 0 u1 0 -5.19165746463552e-06
Rx18 x18 0 1
Fxc18_17 x18 0 Vx17 -1462.84612246587
Cx18 x18 xm18 9.26132475048371e-14
Vx18 xm18 0 0
Gx18_1 x18 0 u1 0 0.00759459599131306
Rx19 x19 0 1
Fxc19_20 x19 0 Vx20 328.769768579133
Cx19 x19 xm19 5.66336887557543e-14
Vx19 xm19 0 0
Gx19_1 x19 0 u1 0 -1.9034828300684e-06
Rx20 x20 0 1
Fxc20_19 x20 0 Vx19 -2278.50862110377
Cx20 x20 xm20 5.66336887557543e-14
Vx20 xm20 0 0
Gx20_1 x20 0 u1 0 0.00433710203843386
Gyc1_1 y1 0 x1 0 1
Gyc1_2 y1 0 x2 0 1
Gyc1_3 y1 0 x3 0 -1
Gyc1_4 y1 0 x4 0 -1
Gyc1_5 y1 0 x5 0 -1
Gyc1_6 y1 0 x6 0 -1
Gyc1_7 y1 0 x7 0 -1
Gyc1_8 y1 0 x8 0 -1
Gyc1_9 y1 0 x9 0 -1
Gyc1_10 y1 0 x10 0 1
Gyc1_11 y1 0 x11 0 1
Gyc1_12 y1 0 x12 0 -1
Gyc1_13 y1 0 x13 0 1
Gyc1_14 y1 0 x14 0 -1
Gyc1_15 y1 0 x15 0 -1
Gyc1_16 y1 0 x16 0 -1
Gyc1_17 y1 0 x17 0 -1
Gyc1_18 y1 0 x18 0 -1
Gyc1_19 y1 0 x19 0 -1
Gyc1_20 y1 0 x20 0 -1
.ENDS
