* Equivalent circuit model for JWS_InductorRed_v2.ckt
.SUBCKT JWS_InductorRed_v2 po1
Vsp1 po1 p1 0
Vsr1 p1 pr1 0
Rp1 pr1 0 50
Ru1 u1 0 50
Fr1 u1 0 Vsr1 -1
Fu1 u1 0 Vsp1 -1
Ry1 y1 0 1
Gy1 p1 0 y1 0 -0.02
Rx1 x1 0 1
Cx1 x1 0 0.018119524928678
Gx1_1 x1 0 u1 0 -2.48050209321686
Rx2 x2 0 1
Cx2 x2 0 0.0462420852993167
Gx2_1 x2 0 u1 0 -3.53224740307816
Rx3 x3 0 1
Fxc3_4 x3 0 Vx4 207.398640746746
Cx3 x3 xm3 0.000177459977133997
Vx3 xm3 0 0
Gx3_1 x3 0 u1 0 -6.29099037658877e-06
Rx4 x4 0 1
Fxc4_3 x4 0 Vx3 -1185.34831840039
Cx4 x4 xm4 0.000177459977133997
Vx4 xm4 0 0
Gx4_1 x4 0 u1 0 0.00745701486396254
Rx5 x5 0 1
Fxc5_6 x5 0 Vx6 404.538373773159
Cx5 x5 xm5 0.000443567499652438
Vx5 xm5 0 0
Gx5_1 x5 0 u1 0 -2.6539583281904e-05
Rx6 x6 0 1
Fxc6_5 x6 0 Vx5 -285.674315648811
Cx6 x6 xm6 0.000443567499652438
Vx6 xm6 0 0
Gx6_1 x6 0 u1 0 0.00758167729166257
Rx7 x7 0 1
Cx7 x7 0 6.23601496088774
Gx7_1 x7 0 u1 0 -2.03850289397003
Gyc1_1 y1 0 x1 0 1
Gyc1_2 y1 0 x2 0 -1
Gyc1_3 y1 0 x3 0 1
Gyc1_4 y1 0 x4 0 -1
Gyc1_5 y1 0 x5 0 1
Gyc1_6 y1 0 x6 0 -1
Gyc1_7 y1 0 x7 0 1
.ENDS
