* Equivalent circuit model for JWS_MixedLoad_v3.ckt
.SUBCKT JWS_MixedLoad_v3 po1
Vsp1 po1 p1 0
Vsr1 p1 pr1 0
Rp1 pr1 0 50
Ru1 u1 0 50
Fr1 u1 0 Vsr1 -1
Fu1 u1 0 Vsp1 -1
Ry1 y1 0 1
Gy1 p1 0 y1 0 -0.02
Rx1 x1 0 1
Cx1 x1 0 8.64470578243862e-12
Gx1_1 x1 0 u1 0 -1.53511965547538
Rx2 x2 0 1
Fxc2_3 x2 0 Vx3 14.2755533077705
Cx2 x2 xm2 1.47644457096936e-12
Vx2 xm2 0 0
Gx2_1 x2 0 u1 0 -0.0284816347070065
Rx3 x3 0 1
Fxc3_2 x3 0 Vx2 -6.09700032467308
Cx3 x3 xm3 1.47644457096936e-12
Vx3 xm3 0 0
Gx3_1 x3 0 u1 0 0.173652536055839
Rx4 x4 0 1
Fxc4_5 x4 0 Vx5 57600.8282085149
Cx4 x4 xm4 7.36226546135046e-16
Vx4 xm4 0 0
Gx4_1 x4 0 u1 0 -7.6022483248364e-09
Rx5 x5 0 1
Fxc5_4 x5 0 Vx4 -8128.75210226842
Cx5 x5 xm5 7.36226546135046e-16
Vx5 xm5 0 0
Gx5_1 x5 0 u1 0 6.17967920524804e-05
Rx6 x6 0 1
Fxc6_7 x6 0 Vx7 51536.8932174199
Cx6 x6 xm6 7.7545696456486e-16
Vx6 xm6 0 0
Gx6_1 x6 0 u1 0 -1.08734732264744e-08
Rx7 x7 0 1
Fxc7_6 x7 0 Vx6 -8283.73149829265
Cx7 x7 xm7 7.75456964564859e-16
Vx7 xm7 0 0
Gx7_1 x7 0 u1 0 9.00729326619874e-05
Rx8 x8 0 1
Fxc8_9 x8 0 Vx9 18645.3851607656
Cx8 x8 xm8 1.69144429889851e-14
Vx8 xm8 0 0
Gx8_1 x8 0 u1 0 -4.17514044985495e-06
Rx9 x9 0 1
Fxc9_8 x9 0 Vx8 -51.9267110859127
Cx9 x9 xm9 1.69144429889851e-14
Vx9 xm9 0 0
Gx9_1 x9 0 u1 0 0.000216801311882726
Rx10 x10 0 1
Fxc10_11 x10 0 Vx11 730.25412135313
Cx10 x10 xm10 1.68365786808145e-13
Vx10 xm10 0 0
Gx10_1 x10 0 u1 0 -0.000464774788536779
Rx11 x11 0 1
Fxc11_10 x11 0 Vx10 -14.9173799531865
Cx11 x11 xm11 1.68365786808145e-13
Vx11 xm11 0 0
Gx11_1 x11 0 u1 0 0.00693322211326506
Rx12 x12 0 1
Fxc12_13 x12 0 Vx13 1107.50465581074
Cx12 x12 xm12 2.08214018407535e-14
Vx12 xm12 0 0
Gx12_1 x12 0 u1 0 -5.43970515054924e-06
Rx13 x13 0 1
Fxc13_12 x13 0 Vx12 -648.961422060721
Cx13 x13 xm13 2.08214018407535e-14
Vx13 xm13 0 0
Gx13_1 x13 0 u1 0 0.00353015879009147
Rx14 x14 0 1
Fxc14_15 x14 0 Vx15 8372.85166951717
Cx14 x14 xm14 1.02910304470458e-14
Vx14 xm14 0 0
Gx14_1 x14 0 u1 0 -1.1370862072317e-06
Rx15 x15 0 1
Fxc15_14 x15 0 Vx14 -411.744978012553
Cx15 x15 xm15 1.02910304470458e-14
Vx15 xm15 0 0
Gx15_1 x15 0 u1 0 0.000468189535394993
Rx16 x16 0 1
Cx16 x16 0 2.28994722979608e-10
Gx16_1 x16 0 u1 0 -2.90593811238065
Rx17 x17 0 1
Fxc17_18 x17 0 Vx18 5098.66572422172
Cx17 x17 xm17 5.33117264892284e-14
Vx17 xm17 0 0
Gx17_1 x17 0 u1 0 -4.52983523619801e-08
Rx18 x18 0 1
Fxc18_17 x18 0 Vx17 -960.453394889496
Cx18 x18 xm18 5.33117264892284e-14
Vx18 xm18 0 0
Gx18_1 x18 0 u1 0 4.35069563089644e-05
Rx19 x19 0 1
Fxc19_20 x19 0 Vx20 5.42809399164623
Cx19 x19 xm19 1.7882319865348e-11
Vx19 xm19 0 0
Gx19_1 x19 0 u1 0 -0.64260650425958
Rx20 x20 0 1
Fxc20_19 x20 0 Vx19 -1.28743405225749
Cx20 x20 xm20 1.7882319865348e-11
Vx20 xm20 0 0
Gx20_1 x20 0 u1 0 0.827313495785932
Rx21 x21 0 1
Fxc21_22 x21 0 Vx22 10556.7284306198
Cx21 x21 xm21 1.80838021682155e-15
Vx21 xm21 0 0
Gx21_1 x21 0 u1 0 -5.18151053505916e-10
Rx22 x22 0 1
Fxc22_21 x22 0 Vx21 -113776.544154347
Cx22 x22 xm22 1.80838021682155e-15
Vx22 xm22 0 0
Gx22_1 x22 0 u1 0 5.89534362178374e-05
Rx23 x23 0 1
Fxc23_24 x23 0 Vx24 17048.6428922445
Cx23 x23 xm23 4.60400202073435e-15
Vx23 xm23 0 0
Gx23_1 x23 0 u1 0 -1.80784452203992e-07
Rx24 x24 0 1
Fxc24_23 x24 0 Vx23 -1267.3240086028
Cx24 x24 xm24 4.60400202073435e-15
Vx24 xm24 0 0
Gx24_1 x24 0 u1 0 0.000229112476660224
Rx25 x25 0 1
Fxc25_26 x25 0 Vx26 581.530173270319
Cx25 x25 xm25 1.76421199618044e-14
Vx25 xm25 0 0
Gx25_1 x25 0 u1 0 -2.7254628077259e-07
Rx26 x26 0 1
Fxc26_25 x26 0 Vx25 -6992.28905717751
Cx26 x26 xm26 1.76421199618044e-14
Vx26 xm26 0 0
Gx26_1 x26 0 u1 0 0.00190572237662061
Rx27 x27 0 1
Fxc27_28 x27 0 Vx28 5971.98398714566
Cx27 x27 xm27 2.55479977751243e-15
Vx27 xm27 0 0
Gx27_1 x27 0 u1 0 -6.84084365201046e-09
Rx28 x28 0 1
Fxc28_27 x28 0 Vx27 -30469.5463813334
Cx28 x28 xm28 2.55479977751243e-15
Vx28 xm28 0 0
Gx28_1 x28 0 u1 0 0.000208437402942383
Rx29 x29 0 1
Fxc29_30 x29 0 Vx30 77.7698128435997
Cx29 x29 xm29 5.46048773523102e-13
Vx29 xm29 0 0
Gx29_1 x29 0 u1 0 -0.00151594257717576
Rx30 x30 0 1
Fxc30_29 x30 0 Vx29 -30.7545776646079
Cx30 x30 xm30 5.46048773523102e-13
Vx30 xm30 0 0
Gx30_1 x30 0 u1 0 0.0466221737248377
Rx31 x31 0 1
Fxc31_32 x31 0 Vx32 614.336845196194
Cx31 x31 xm31 1.46477096533141e-14
Vx31 xm31 0 0
Gx31_1 x31 0 u1 0 -4.90571152420862e-07
Rx32 x32 0 1
Fxc32_31 x32 0 Vx31 -4633.6579328877
Cx32 x32 xm32 1.46477096533141e-14
Vx32 xm32 0 0
Gx32_1 x32 0 u1 0 0.00227313891206079
Rx33 x33 0 1
Fxc33_34 x33 0 Vx34 438.455282604189
Cx33 x33 xm33 4.20876591287536e-14
Vx33 xm33 0 0
Gx33_1 x33 0 u1 0 -6.9671282538441e-06
Rx34 x34 0 1
Fxc34_33 x34 0 Vx33 -804.307146043073
Cx34 x34 xm34 4.20876591287536e-14
Vx34 xm34 0 0
Gx34_1 x34 0 u1 0 0.00560371104196541
Gyc1_1 y1 0 x1 0 1
Gyc1_2 y1 0 x2 0 -1
Gyc1_3 y1 0 x3 0 -1
Gyc1_4 y1 0 x4 0 -1
Gyc1_5 y1 0 x5 0 1
Gyc1_6 y1 0 x6 0 -1
Gyc1_7 y1 0 x7 0 1
Gyc1_8 y1 0 x8 0 -1
Gyc1_9 y1 0 x9 0 1
Gyc1_10 y1 0 x10 0 -1
Gyc1_11 y1 0 x11 0 1
Gyc1_12 y1 0 x12 0 1
Gyc1_13 y1 0 x13 0 1
Gyc1_14 y1 0 x14 0 -1
Gyc1_15 y1 0 x15 0 1
Gyc1_16 y1 0 x16 0 -1
Gyc1_17 y1 0 x17 0 -1
Gyc1_18 y1 0 x18 0 1
Gyc1_19 y1 0 x19 0 -1
Gyc1_20 y1 0 x20 0 -1
Gyc1_21 y1 0 x21 0 1
Gyc1_22 y1 0 x22 0 1
Gyc1_23 y1 0 x23 0 -1
Gyc1_24 y1 0 x24 0 -1
Gyc1_25 y1 0 x25 0 -1
Gyc1_26 y1 0 x26 0 -1
Gyc1_27 y1 0 x27 0 -1
Gyc1_28 y1 0 x28 0 -1
Gyc1_29 y1 0 x29 0 -1
Gyc1_30 y1 0 x30 0 -1
Gyc1_31 y1 0 x31 0 -1
Gyc1_32 y1 0 x32 0 -1
Gyc1_33 y1 0 x33 0 -1
Gyc1_34 y1 0 x34 0 -1
.ENDS
