* Equivalent circuit model for kimball_10MHzto3p3GHz_R50.ckt
.SUBCKT kimball_10MHzto3p3GHz_R50 po1
Vsp1 po1 p1 0
Eu1 u1 um1 p1 0 1
Hu1 um1 0 Vsp1 50
Ru1 u1 0 1
Rx1 x1 0 1
Cx1 x1 xm1 2.66711857033722e-11
Vx1 xm1 0 0
Fxc1_2 x1 0 Vx2 0.426471344009162
Gx1_1 x1 0 u1 0 -0.417210152499289
Rx2 x2 0 1
Cx2 x2 xm2 2.66711857033722e-11
Vx2 xm2 0 0
Fxc2_1 x2 0 Vx1 -3.0073443607057
Gx2_1 x2 0 u1 0 1.2546945993479
Rx3 x3 0 1
Cx3 x3 xm3 5.56070623565171e-12
Vx3 xm3 0 0
Fxc3_4 x3 0 Vx4 6.75999740840829
Gx3_1 x3 0 u1 0 -0.037767671988619
Rx4 x4 0 1
Cx4 x4 xm4 5.56070623565171e-12
Vx4 xm4 0 0
Fxc4_3 x4 0 Vx3 -10.7671658026464
Gx4_1 x4 0 u1 0 0.406650786281426
Rx5 x5 0 1
Cx5 x5 xm5 4.42300002509665e-14
Vx5 xm5 0 0
Fxc5_6 x5 0 Vx6 1312.96417088542
Gx5_1 x5 0 u1 0 -2.00693860567888e-06
Rx6 x6 0 1
Cx6 x6 xm6 4.42300002509665e-14
Vx6 xm6 0 0
Fxc6_5 x6 0 Vx5 -1126.13956510721
Gx6_1 x6 0 u1 0 0.00226009296859609
Rx7 x7 0 1
Cx7 x7 xm7 6.03253163057338e-10
Vx7 xm7 0 0
Gx7_1 x7 0 u1 0 -2.23099332608783
Ry1 y1 0 1
Gyc1_1 y1 0 x1 0 1
Gyc1_2 y1 0 x2 0 -1
Gyc1_3 y1 0 x3 0 -1
Gyc1_4 y1 0 x4 0 1
Gyc1_5 y1 0 x5 0 1
Gyc1_6 y1 0 x6 0 1
Gyc1_7 y1 0 x7 0 -1
Ey1 p1 0 y1 ym1 1
Hy1 ym1 0 Vsp1 -50
.ENDS
