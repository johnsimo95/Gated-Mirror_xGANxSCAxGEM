* Equivalent circuit model for JWS_InductorRed_v6.ckt
.SUBCKT JWS_InductorRed_v6 po1
Vsp1 po1 p1 0
Vsr1 p1 pr1 0
Rp1 pr1 0 50
Ru1 u1 0 50
Fr1 u1 0 Vsr1 -1
Fu1 u1 0 Vsp1 -1
Ry1 y1 0 1
Gy1 p1 0 y1 0 -0.02
Rx1 x1 0 1
Fxc1_2 x1 0 Vx2 1.35233127278082
Cx1 x1 xm1 0.00699985480109497
Vx1 xm1 0 0
Gx1_1 x1 0 u1 0 -0.675796516388234
Rx2 x2 0 1
Fxc2_1 x2 0 Vx1 -1.00698059719778
Cx2 x2 xm2 0.00699985480109497
Vx2 xm2 0 0
Gx2_1 x2 0 u1 0 0.680513979656805
Rx3 x3 0 1
Fxc3_4 x3 0 Vx4 532.367812664324
Cx3 x3 xm3 0.000100763821370372
Vx3 xm3 0 0
Gx3_1 x3 0 u1 0 -0.000106386911571397
Rx4 x4 0 1
Fxc4_3 x4 0 Vx3 -47.3623505456546
Cx4 x4 xm4 0.000100763821370372
Vx4 xm4 0 0
Gx4_1 x4 0 u1 0 0.00503873419931406
Rx5 x5 0 1
Fxc5_6 x5 0 Vx6 6303.70087058227
Cx5 x5 xm5 3.45266372683876e-06
Vx5 xm5 0 0
Gx5_1 x5 0 u1 0 -1.26255625339998e-07
Rx6 x6 0 1
Fxc6_5 x6 0 Vx5 -3967.67362295263
Cx6 x6 xm6 3.45266372683877e-06
Vx6 xm6 0 0
Gx6_1 x6 0 u1 0 0.000500941114410898
Rx7 x7 0 1
Fxc7_8 x7 0 Vx8 738.456864533614
Cx7 x7 xm7 6.3245698301244e-05
Vx7 xm7 0 0
Gx7_1 x7 0 u1 0 -5.33601329095001e-05
Rx8 x8 0 1
Fxc8_7 x8 0 Vx7 -104.213495994539
Cx8 x8 xm8 6.3245698301244e-05
Vx8 xm8 0 0
Gx8_1 x8 0 u1 0 0.00556084599723227
Rx9 x9 0 1
Fxc9_10 x9 0 Vx10 2306.53041673434
Cx9 x9 xm9 6.79328432793681e-06
Vx9 xm9 0 0
Gx9_1 x9 0 u1 0 -4.21198302199632e-07
Rx10 x10 0 1
Fxc10_9 x10 0 Vx9 -2924.36622091829
Cx10 x10 xm10 6.79328432793681e-06
Vx10 xm10 0 0
Gx10_1 x10 0 u1 0 0.00123173808726074
Rx11 x11 0 1
Fxc11_12 x11 0 Vx12 2840.13554850218
Cx11 x11 xm11 5.42942223317773e-05
Vx11 xm11 0 0
Gx11_1 x11 0 u1 0 -3.56363186967412e-05
Rx12 x12 0 1
Fxc12_11 x12 0 Vx11 -40.1977701236042
Cx12 x12 xm12 5.42942223317773e-05
Vx12 xm12 0 0
Gx12_1 x12 0 u1 0 0.0014325005470231
Rx13 x13 0 1
Fxc13_14 x13 0 Vx14 411.316004608491
Cx13 x13 xm13 0.000150605509895977
Vx13 xm13 0 0
Gx13_1 x13 0 u1 0 -0.000213633334438348
Rx14 x14 0 1
Fxc14_13 x14 0 Vx13 -44.5476486636099
Cx14 x14 xm14 0.000150605509895977
Vx14 xm14 0 0
Gx14_1 x14 0 u1 0 0.00951686272539501
Rx15 x15 0 1
Fxc15_16 x15 0 Vx16 49263.111806473
Cx15 x15 xm15 3.40517599500512e-06
Vx15 xm15 0 0
Gx15_1 x15 0 u1 0 -9.94531123401774e-08
Rx16 x16 0 1
Fxc16_15 x16 0 Vx15 -789.777680542131
Cx16 x16 xm16 3.40517599500512e-06
Vx16 xm16 0 0
Gx16_1 x16 0 u1 0 7.85458483867213e-05
Rx17 x17 0 1
Cx17 x17 0 0.0525968036428866
Gx17_1 x17 0 u1 0 -2.47462910655772
Rx18 x18 0 1
Fxc18_19 x18 0 Vx19 628.47384793395
Cx18 x18 xm18 7.90266093469789e-05
Vx18 xm18 0 0
Gx18_1 x18 0 u1 0 -4.66110054961111e-05
Rx19 x19 0 1
Fxc19_18 x19 0 Vx18 -128.551740640618
Cx19 x19 xm19 7.90266093469789e-05
Vx19 xm19 0 0
Gx19_1 x19 0 u1 0 0.00599192588953448
Rx20 x20 0 1
Fxc20_21 x20 0 Vx21 17387.5803105237
Cx20 x20 xm20 1.62645751439864e-05
Vx20 xm20 0 0
Gx20_1 x20 0 u1 0 -2.04720033949162e-06
Rx21 x21 0 1
Fxc21_20 x21 0 Vx20 -113.88435170192
Cx21 x21 xm21 1.62645751439864e-05
Vx21 xm21 0 0
Gx21_1 x21 0 u1 0 0.000233144083466954
Rx22 x22 0 1
Fxc22_23 x22 0 Vx23 350.818300586562
Cx22 x22 xm22 0.0002070143232839
Vx22 xm22 0 0
Gx22_1 x22 0 u1 0 -0.000273487642402542
Rx23 x23 0 1
Fxc23_22 x23 0 Vx22 -40.5328906510395
Cx23 x23 xm23 0.000207014323283901
Vx23 xm23 0 0
Gx23_1 x23 0 u1 0 0.0110852447039128
Rx24 x24 0 1
Fxc24_25 x24 0 Vx25 26596.5575931445
Cx24 x24 xm24 2.34051275503381e-06
Vx24 xm24 0 0
Gx24_1 x24 0 u1 0 -2.91778131711961e-08
Rx25 x25 0 1
Fxc25_24 x25 0 Vx24 -4944.98966267492
Cx25 x25 xm25 2.34051275503381e-06
Vx25 xm25 0 0
Gx25_1 x25 0 u1 0 0.000144283984511025
Rx26 x26 0 1
Fxc26_27 x26 0 Vx27 7171.8446519837
Cx26 x26 xm26 1.01830191819747e-05
Vx26 xm26 0 0
Gx26_1 x26 0 u1 0 -5.21712548206203e-07
Rx27 x27 0 1
Fxc27_26 x27 0 Vx26 -994.401002678934
Cx27 x27 xm27 1.01830191819747e-05
Vx27 xm27 0 0
Gx27_1 x27 0 u1 0 0.000518791481046429
Rx28 x28 0 1
Cx28 x28 0 6.19795566853536
Gx28_1 x28 0 u1 0 -2.03540901112705
Rx29 x29 0 1
Fxc29_30 x29 0 Vx30 400.479978643746
Cx29 x29 xm29 0.000444944006147345
Vx29 xm29 0 0
Gx29_1 x29 0 u1 0 -2.65066745220706e-05
Rx30 x30 0 1
Fxc30_29 x30 0 Vx29 -286.783458443473
Cx30 x30 xm30 0.000444944006147345
Vx30 xm30 0 0
Gx30_1 x30 0 u1 0 0.00760167579127491
Rx31 x31 0 1
Fxc31_32 x31 0 Vx32 207.548812431025
Cx31 x31 xm31 0.000177462968015681
Vx31 xm31 0 0
Gx31_1 x31 0 u1 0 -6.27748545270282e-06
Rx32 x32 0 1
Fxc32_31 x32 0 Vx31 -1184.44589894556
Cx32 x32 xm32 0.000177462968015681
Vx32 xm32 0 0
Gx32_1 x32 0 u1 0 0.00743534190014425
Rx33 x33 0 1
Fxc33_34 x33 0 Vx34 31858.0917834618
Cx33 x33 xm33 1.22288686325781e-06
Vx33 xm33 0 0
Gx33_1 x33 0 u1 0 -3.18542166963733e-09
Rx34 x34 0 1
Fxc34_33 x34 0 Vx33 -18392.8408192811
Cx34 x34 xm34 1.22288686325781e-06
Vx34 xm34 0 0
Gx34_1 x34 0 u1 0 5.85889537119279e-05
Rx35 x35 0 1
Fxc35_36 x35 0 Vx36 408.223073797884
Cx35 x35 xm35 9.22840667656988e-05
Vx35 xm35 0 0
Gx35_1 x35 0 u1 0 -2.56000982655997e-05
Rx36 x36 0 1
Fxc36_35 x36 0 Vx35 -293.484880047035
Cx36 x36 xm36 9.22840667656988e-05
Vx36 xm36 0 0
Gx36_1 x36 0 u1 0 0.00751324176867184
Rx37 x37 0 1
Fxc37_38 x37 0 Vx38 4314.76898313907
Cx37 x37 xm37 8.19921701916302e-06
Vx37 xm37 0 0
Gx37_1 x37 0 u1 0 -1.6622347883535e-07
Rx38 x38 0 1
Fxc38_37 x38 0 Vx37 -4111.96936104881
Cx38 x38 xm38 8.19921701916302e-06
Vx38 xm38 0 0
Gx38_1 x38 0 u1 0 0.000683505852057903
Rx39 x39 0 1
Fxc39_40 x39 0 Vx40 1977.02495881025
Cx39 x39 xm39 1.45799045367297e-05
Vx39 xm39 0 0
Gx39_1 x39 0 u1 0 -3.7778516870885e-07
Rx40 x40 0 1
Fxc40_39 x40 0 Vx39 -3324.75024958692
Cx40 x40 xm40 1.45799045367297e-05
Vx40 xm40 0 0
Gx40_1 x40 0 u1 0 0.00125604133395498
Rx41 x41 0 1
Fxc41_42 x41 0 Vx42 293.397710510842
Cx41 x41 xm41 1.04392969223032e-05
Vx41 xm41 0 0
Gx41_1 x41 0 u1 0 -7.81893114818686e-09
Rx42 x42 0 1
Fxc42_41 x42 0 Vx41 -112343.096952249
Cx42 x42 xm42 1.04392969223032e-05
Vx42 xm42 0 0
Gx42_1 x42 0 u1 0 0.00087840294004372
Rx43 x43 0 1
Fxc43_44 x43 0 Vx44 173.100470195996
Cx43 x43 xm43 9.19239040861538e-05
Vx43 xm43 0 0
Gx43_1 x43 0 u1 0 -5.1333222420833e-06
Rx44 x44 0 1
Fxc44_43 x44 0 Vx43 -1468.26544339181
Cx44 x44 xm44 9.19239040861538e-05
Vx44 xm44 0 0
Gx44_1 x44 0 u1 0 0.00753707965784547
Rx45 x45 0 1
Fxc45_46 x45 0 Vx46 764.257205268387
Cx45 x45 xm45 0.000136119595064061
Vx45 xm45 0 0
Gx45_1 x45 0 u1 0 -5.23192082740176e-06
Rx46 x46 0 1
Fxc46_45 x46 0 Vx45 -169.848789574195
Cx46 x46 xm46 0.000136119595064061
Vx46 xm46 0 0
Gx46_1 x46 0 u1 0 0.000888635419682211
Rx47 x47 0 1
Fxc47_48 x47 0 Vx48 494.265313449122
Cx47 x47 xm47 6.81122506914562e-05
Vx47 xm47 0 0
Gx47_1 x47 0 u1 0 -4.67645965081204e-06
Rx48 x48 0 1
Fxc48_47 x48 0 Vx47 -1047.55561635742
Cx48 x48 xm48 6.81122506914562e-05
Vx48 xm48 0 0
Gx48_1 x48 0 u1 0 0.00489885157187702
Gyc1_1 y1 0 x1 0 1
Gyc1_2 y1 0 x2 0 -1
Gyc1_3 y1 0 x3 0 -1
Gyc1_4 y1 0 x4 0 -1
Gyc1_5 y1 0 x5 0 -1
Gyc1_6 y1 0 x6 0 -1
Gyc1_7 y1 0 x7 0 -1
Gyc1_8 y1 0 x8 0 -1
Gyc1_9 y1 0 x9 0 -1
Gyc1_10 y1 0 x10 0 1
Gyc1_11 y1 0 x11 0 -1
Gyc1_12 y1 0 x12 0 -1
Gyc1_13 y1 0 x13 0 -1
Gyc1_14 y1 0 x14 0 -1
Gyc1_15 y1 0 x15 0 -1
Gyc1_16 y1 0 x16 0 -1
Gyc1_17 y1 0 x17 0 -1
Gyc1_18 y1 0 x18 0 -1
Gyc1_19 y1 0 x19 0 -1
Gyc1_20 y1 0 x20 0 -1
Gyc1_21 y1 0 x21 0 -1
Gyc1_22 y1 0 x22 0 -1
Gyc1_23 y1 0 x23 0 -1
Gyc1_24 y1 0 x24 0 -1
Gyc1_25 y1 0 x25 0 -1
Gyc1_26 y1 0 x26 0 -1
Gyc1_27 y1 0 x27 0 -1
Gyc1_28 y1 0 x28 0 1
Gyc1_29 y1 0 x29 0 1
Gyc1_30 y1 0 x30 0 -1
Gyc1_31 y1 0 x31 0 1
Gyc1_32 y1 0 x32 0 -1
Gyc1_33 y1 0 x33 0 -1
Gyc1_34 y1 0 x34 0 -1
Gyc1_35 y1 0 x35 0 -1
Gyc1_36 y1 0 x36 0 -1
Gyc1_37 y1 0 x37 0 -1
Gyc1_38 y1 0 x38 0 -1
Gyc1_39 y1 0 x39 0 -1
Gyc1_40 y1 0 x40 0 -1
Gyc1_41 y1 0 x41 0 -1
Gyc1_42 y1 0 x42 0 -1
Gyc1_43 y1 0 x43 0 -1
Gyc1_44 y1 0 x44 0 -1
Gyc1_45 y1 0 x45 0 1
Gyc1_46 y1 0 x46 0 1
Gyc1_47 y1 0 x47 0 -1
Gyc1_48 y1 0 x48 0 -1
.ENDS
